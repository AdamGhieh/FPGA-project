library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity i_cache is
port (
    address_input : in std_logic_vector(31 downto 0);
    data_output : out std_logic_vector(31 downto 0)
);
end i_cache;

architecture behav of i_cache is
begin
    process (address_input)
    begin
        case address_input is
		
            when x"00000000" => data_output <= x"00000113"; -- addi x2,x0,0
            when x"00000004" => data_output <= x"00500193"; -- addi x3,x0,5
            when x"00000008" => data_output <= x"00000217"; -- auipc x4, 0
            when x"0000000C" => data_output <= x"00316663"; -- loop: bltu x2, x3, store
            when x"00000010" => data_output <= x"0180026F"; -- jal x4, function
            when x"00000014" => data_output <= x"00000063"; -- done: beq x0, x0, done
            when x"00000018" => data_output <= x"02410823"; -- store: sb x4, 0x30(x2)
            when x"0000001C" => data_output <= x"00110113"; -- addi x2, x2, 1
            when x"00000020" => data_output <= x"00121213"; -- slli x4, x4, 1
            when x"00000024" => data_output <= x"FE9FF06F"; -- jal x0, loop
            when x"00000028" => data_output <= x"03404283"; -- funtion: lbu x5, 0x34(x0)
            when x"0000002C" => data_output <= x"0002A313"; -- slti x6, x5, 0
            when x"00000030" => data_output <= x"03400283"; -- lb, x5, 0x34(x0) 
            when x"00000034" => data_output <= x"0002A393"; -- slti x7, x5, 0
            when x"00000038" => data_output <= x"00730A63"; -- beq x6, x7, error
            when x"0000003C" => data_output <= x"4012D293"; -- srai x5, x5, 1
            when x"00000040" => data_output <= x"FbF00313"; -- addi x6, x0, -65
            when x"00000044" => data_output <= x"00535463"; -- bge x6, x5, error
            when x"00000048" => data_output <= x"00020067"; -- jalr x0, 0(x4)
            when x"0000004C" => data_output <= x"00000063"; -- error: beq x0, x0, error
            when others => data_output <= x"00000000"; -- don't care
        end case;
    end process;
end behav;
